module not1(input i1, output o1);
  assign o1 = !i1;
endmodule
